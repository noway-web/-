`timescale 1ns / 1ps

module testbench();

// Регистры и проводники для тестирования
reg [5:0] args;              // Регистр для хранения аргументов
reg clk;                     // Регистр для симуляции тактового сигнала
wire res1, res2;                    // Выходной проводник (результат)
reg [0:31] reference_reg, error_reg1, error_reg2;    // Регистр для хранения эталонных данных, регистр для хранения ошибок

initial
begin
    reference_reg = 32'hD5BA8AE9;  // Инициализация эталонного регистра
    args = 5'b00000;             // Инициализация аргументов
    clk = 0;                     // Инициализация симуляции тактового сигнала
    error_reg1 = 0;               // Инициализация регистра ошибок
    error_reg2 = 0;               // Инициализация регистра ошибок
end

// Генерация тактового сигнала с периодом 10 временных единиц
always #10 clk = ~clk;

// Обработка на каждом положительном фронте тактового сигнала
always @(posedge clk)
begin
    error_reg1[args] = res1 ~^ reference_reg[args];  // Вычисление ошибки для текущего аргумента
    error_reg2[args] = res2 ~^ reference_reg[args];
    args = args + 1;                              // Увеличение аргумента на 1
    if(args == 6'd33)
        $finish;                                   // Завершение симуляции после обработки всех аргументов
end      
sdnf mod1 (.in(args[4:0]), .f(res1));          // Вызов модуля "main_sdnf" с текущим аргументом
mdnf mod2 (.in(args[4:0]), .f(res2));  
endmodule
