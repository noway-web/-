`timescale 1ns / 1ps

module sdnf (
    input wire [4:0] in,   // Входной сигнал in состоит из 5 бит
    output wire f          // Выходной сигнал f
);

assign f = (~in[4] & ~in[3] & ~in[2] & ~in[1] & ~in[0]) // K1: { 0, 0, 0, 0, 0 } — ¬x1¬x2¬x3¬x4¬x5
           || (~in[4] & ~in[3] & ~in[2] & ~in[1] & in[0]) // K2: { 0, 0, 0, 0, 1 } — ¬x1¬x2¬x3¬x4x5
           || (~in[4] & ~in[3] & ~in[2] & in[1] & in[0]) // K3: { 0, 0, 0, 1, 1 } — ¬x1¬x2¬x3x4x5
           || (~in[4] & ~in[3] & in[2] & ~in[1] & in[0]) // K4: { 0, 0, 1, 0, 1 } — ¬x1¬x2x3¬x4x5
           || (~in[4] & ~in[3] & in[2] & in[1] & in[0]) // K5: { 0, 0, 1, 1, 1 } — ¬x1¬x2x3x4x5
           || (~in[4] & in[3] & ~in[2] & ~in[1] & ~in[0]) // K6: { 0, 1, 0, 0, 0 } — ¬x1x2¬x3¬x4¬x5
           || (~in[4] & in[3] & ~in[2] & ~in[1] & in[0]) // K7: { 0, 1, 0, 1, 0 } — ¬x1x2¬x3x4¬x5
           || (~in[4] & in[3] & ~in[2] & in[1] & in[0]) // K8: { 0, 1, 0, 1, 1 } — ¬x1x2¬x3x4x5
           || (~in[4] & in[3] & in[2] & ~in[1] & ~in[0]) // K9: { 0, 1, 1, 0, 0 } — ¬x1x2x3¬x4¬x5
           || (~in[4] & in[3] & in[2] & in[1] & ~in[0]) // K10: { 0, 1, 1, 1, 0 } — ¬x1x2x3x4¬x5
           || (in[4] & ~in[3] & ~in[2] & ~in[1] & ~in[0]) // K11: { 1, 0, 0, 0, 0 } — x1¬x2¬x3¬x4¬x5
           || (in[4] & ~in[3] & in[2] & ~in[1] & ~in[0]) // K12: { 1, 0, 1, 0, 0 } — x1¬x2x3¬x4¬x5
           || (in[4] & ~in[3] & in[2] & in[1] & ~in[0]) // K13: { 1, 0, 1, 1, 0 } — x1¬x2x3x4¬x5
           || (in[4] & in[3] & ~in[2] & ~in[1] & ~in[0]) // K14: { 1, 1, 0, 0, 0 } — x1x2¬x3¬x4¬x5
           || (in[4] & in[3] & ~in[2] & ~in[1] & in[0]) // K15: { 1, 1, 0, 0, 1 } — x1x2¬x3¬x4x5
           || (in[4] & in[3] & ~in[2] & in[1] & ~in[0]) // K16: { 1, 1, 0, 1, 0 } — x1x2¬x3x4¬x5
           || (in[4] & in[3] & in[2] & ~in[1] & ~in[0]) // K17: { 1, 1, 1, 0, 0 } — x1x2x3¬x4¬x5
           || (in[4] & in[3] & in[2] & in[1] & in[0]); // K18: { 1, 1, 1, 1, 1 } — x1x2x3x4x5
          
endmodule

module mdnf (
    input wire [4:0] in,   // Входной сигнал in состоит из 5 бит
    output wire f          // Выходной сигнал f
);

   assign f = (~in[4] & in[3] & ~in[0]) ||     // ¬x1x2¬x5
               (in[3] & ~in[2] & ~in[0]) ||    // x2¬x3¬x5
               (~in[4] & ~in[3] & in[0]) ||    // ¬x1¬x2x5
               (in[4] & in[3] & ~in[2] & ~in[1]) || // x1x2¬x3¬x4
               (in[4] & ~in[3] & in[2] & ~in[0]) || // x1¬x2x3¬x5
               (in[4] & in[3] & in[2] & in[1] & in[0]) || // x1x2x3x4x5
               (in[4] & ~in[1] & ~in[0]) || // x1¬x4¬x5
               (~in[2] & ~in[1] & ~in[0]) || // ¬x3¬x4¬x5
               (~in[4] & ~in[3] & ~in[2] & in[1]); // ¬x1x2¬x3x4
endmodule
